----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 06/15/2023 05:20:51 PM
-- Design Name: 
-- Module Name: trigger_update - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity trigger_update is
    generic ( CNT_BIT : positive := 16);
    port ( 
        -- >>> OUTPUT >>>
        update_o : out std_logic; -- update trigger generated by the comparator
        -- <<< OUTPUT <<<
        -- >>> INPUT >>>
        max_i :  in std_logic_vector (CNT_BIT-1 downto 0);
        counter_i :  in std_logic_vector (CNT_BIT-1 downto 0);
        peak_i : in std_logic := '0';
        valley_i : in std_logic := '0';
        sawtri_i : in std_logic := '0'
        -- <<< INPUT <<<
        );
end trigger_update;

architecture Behavioral of trigger_update is
    signal maxtrig_s : std_logic;
    signal zerotrig_s : std_logic;
    signal sawtrig_s : std_logic;
    signal tritrig_s : std_logic;
begin
    -- >>> TRIGGER COMPARATORS >>>
    COMPARATOR_MAX : process(counter_i, max_i)
    begin
        if unsigned(counter_i) = unsigned(max_i) then
            maxtrig_s <= '1';
        else
            maxtrig_s <= '0';
        end if;
    end process;
    COMPARATOR_ZERO : process(counter_i)
    begin
        if unsigned(counter_i) = 0 then
            zerotrig_s <= '1';
        else
            zerotrig_s <= '0';
        end if;
    end process;
    -- >>> TRIGGER COMPARATORS >>>
    
    -- >>> TRIGGER SELECTOR >>>
    sawtrig_s <= maxtrig_s;
    tritrig_s <= (maxtrig_s and peak_i) or (zerotrig_s and valley_i);
    
    SAWTRI_TRIGGER : process(sawtri_i, sawtrig_s, tritrig_s)
    begin
        case sawtri_i is
        when '0' => 
            update_o <= sawtrig_s;
        when others =>
            update_o <= tritrig_s;
        end case;
    end process;
    -- >>> TRIGGER SELECTOR >>>
    
end Behavioral;
