----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 06/15/2023 02:16:36 PM
-- Design Name: 
-- Module Name: trigger_generator - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;


entity trigger_generator is
    generic ( CNT_BIT : positive := 16; SEL_BIT : positive := 2);
    port ( 
        -- >>> OUTPUT >>>
        trig_o : out std_logic; -- trigger generated by the comparator
        -- <<< OUTPUT <<<
        -- >>> INPUT >>>
        zero_i : in std_logic_vector (CNT_BIT-1 downto 0);
        first_i : in std_logic_vector (CNT_BIT-1 downto 0);
        second_i : in std_logic_vector (CNT_BIT-1 downto 0);
        third_i :  in std_logic_vector (CNT_BIT-1 downto 0);
        counter_i :  in std_logic_vector (CNT_BIT-1 downto 0);
        sel_i : in std_logic_vector(SEL_BIT-1 downto 0) := (others => '0') -- input value selector | 00=zero | 01=first | etc.
        -- <<< INPUT <<<
        );
end trigger_generator;

architecture Behavioral of trigger_generator is
    type array_mux_t is array (0 to 2**SEL_BIT-1) of std_logic_vector(CNT_BIT-1 downto 0);
    signal mux_a  : array_mux_t;
    signal muxed_s : unsigned(CNT_BIT-1 downto 0);
begin
    -- >>> MULTIPLEXED SELECTOR >>>
    mux_a(0) <= zero_i;
    mux_a(1) <= first_i;
    mux_a(2) <= second_i;
    mux_a(3) <= third_i;
    muxed_s <= unsigned(mux_a(to_integer(unsigned(sel_i))));
    -- <<< MULTIPLEXED SELECTOR <<<
    
    -- >>> TRIGGER COMPARATOR >>>
    COMPARATOR_LOGIC : process(counter_i, muxed_s)
    begin
        if muxed_s = unsigned(counter_i) then
            trig_o <= '1';
        else
            trig_o <= '0';
        end if;
    end process;
    -- <<< TRIGGER COMPARATOR <<<

end Behavioral;
